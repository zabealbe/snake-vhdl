library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sheet_rom is
generic (
    addr_width: integer := 19456;
    data_width: integer := 12
);
port (
    index: in integer range 0 to addr_width - 1;
    data: out std_logic_vector(data_width - 1 downto 0)
);
constant rom_size: integer := 19456;
attribute size: integer;
attribute size of sheet_rom : entity is rom_size;

constant rom_width: integer := 608;
attribute width: integer;
attribute width of sheet_rom : entity is rom_width;

constant rom_height: integer := 32;
attribute height: integer;
attribute height of sheet_rom : entity is rom_height;
end sheet_rom;

architecture Behavioral of sheet_rom is
    type rom_type is array (0 to addr_width - 1) of std_logic_vector(data_width - 1 downto 0);
    signal rom: rom_type := ("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","100001000000","100001000000","100001000000","100001000000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","100001000000","100001000000","100001000000","100001000000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","100001000000","100001000000","100001000000","100001000000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","100001000000","100001000000","100001000000","100001000000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001101100100","001101100100","001101100100","001101100100","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001101100100","001101100100","001101100100","001101100100","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001101100100","001101100100","001101100100","001101100100","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001101100100","001101100100","001101100100","001101100100","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","100001000000","100001000000","100001000000","100001000000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","111111111111","111111111111","111111111111","111111111111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","011111101001","011111101001","011111101001","011111101001","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","111001010000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","111110100000","111110100000","111110100000","111110100000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","100001000000","111110100000","111110100000","111110100000","111110100000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","101000110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","110001110000","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","001000001011","001000001011","001000001011","001000001011","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","010001101111","011010101111","011010101111","011010101111","011010101111","010001101111","010001101111","010001101111","010001101111","001000001011","001000001011","001000001011","001000001011","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111","010110100111");
begin
    data <= rom(index);
end Behavioral; 