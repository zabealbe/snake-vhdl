library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.graphics_pkg.all;

entity tileset_rom is
port (
    tile_index: in integer range 0 to 59 - 1;
    tile_offx: in t_tile_offx;
    tile_offy: in t_tile_offy;
    data: out std_logic_vector(12 - 1 downto 0)
);
end tileset_rom;

architecture Behavioral of tileset_rom is
    type t_rom0 is array (0 to 8 - 1)  of std_logic_vector(12 - 1 downto 0);
    type t_rom1 is array (0 to 8 - 1) of t_rom0;
    type t_rom  is array (0 to 59 - 1) of t_rom1;
    signal rom: t_rom := (
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "000000000000", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "111111111111", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "000000000000", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "000000000000", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "111111111111", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "111111111111", "000000000000", "000000000000"), 
		("000000000000", "000000000000", "111111111111", "111111111111", "111111111111", "000000000000", "000000000000", "000000000000")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "011111101001", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "011111101001", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "001101100100", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "011111101001", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "100001000000", "100001000000", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "100001000000", "100001000000", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "101000110000", "100001000000", "101000110000", "101000110000", "010110100111", "010110100111"), 
		("010110100111", "101000110000", "111001010000", "111001010000", "111001010000", "111001010000", "101000110000", "010110100111"), 
		("010110100111", "101000110000", "111001010000", "111001010000", "111001010000", "111001010000", "101000110000", "010110100111"), 
		("010110100111", "101000110000", "111001010000", "111001010000", "111001010000", "111001010000", "101000110000", "010110100111"), 
		("010110100111", "010110100111", "101000110000", "101000110000", "101000110000", "101000110000", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("110001110000", "110001110000", "110001110000", "110001110000", "110001110000", "110001110000", "110001110000", "110001110000"), 
		("110001110000", "111110100000", "100001000000", "100001000000", "100001000000", "100001000000", "111110100000", "110001110000"), 
		("110001110000", "100001000000", "110001110000", "100001000000", "100001000000", "110001110000", "100001000000", "110001110000"), 
		("110001110000", "100001000000", "100001000000", "110001110000", "100001000000", "100001000000", "100001000000", "110001110000"), 
		("110001110000", "100001000000", "100001000000", "100001000000", "110001110000", "100001000000", "100001000000", "110001110000"), 
		("110001110000", "100001000000", "110001110000", "100001000000", "100001000000", "110001110000", "100001000000", "110001110000"), 
		("110001110000", "111110100000", "100001000000", "100001000000", "100001000000", "100001000000", "111110100000", "110001110000"), 
		("110001110000", "110001110000", "110001110000", "110001110000", "110001110000", "110001110000", "110001110000", "110001110000")
	),
	(
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "000000010000", "010001101111", "010001101111", "000000010000", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "000000010000", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "011010101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "000000010000", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "000000010000", "010001101111", "010001101111", "000000010000", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111")
	),
	(
		("010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "000000010000", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("011010101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "000000010000", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111", "011010101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "011010101111", "010001101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("011010101111", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111")
	),
	(
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "011010101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010001101111", "011010101111", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("011010101111", "010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("010110100111", "010110100111", "001000001011", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111", "011010101111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111"), 
		("010110100111", "010110100111", "001000001011", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "001000001011", "010001101111", "010001101111", "001000001011", "010110100111", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "001000001011", "010110100111", "010110100111"), 
		("010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("011010101111", "010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "001000001011", "001000001011", "010110100111", "010110100111"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("010001101111", "011010101111", "010001101111", "011010101111", "010001101111", "011010101111", "010001101111", "011010101111"), 
		("011010101111", "010001101111", "011010101111", "010001101111", "011010101111", "010001101111", "011010101111", "010001101111"), 
		("010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111", "010001101111"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "001000001011", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "000000010000", "010001101111", "010001101111", "000000010000", "010001101111", "001000001011"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("001000001011", "101000110000", "111111111111", "111001010000", "111001010000", "111111111111", "101000110000", "001000001011"), 
		("010110100111", "101000110000", "111001010000", "111001010000", "111001010000", "111001010000", "101000110000", "010110100111"), 
		("010110100111", "010110100111", "101000110000", "101000110000", "101000110000", "101000110000", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "100001000000", "001000001011", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "010110100111", "101000110000", "111111111111", "001000001011", "000000010000", "010001101111", "010001101111"), 
		("010110100111", "101000110000", "111001010000", "111001010000", "001000001011", "010001101111", "010001101111", "011010101111"), 
		("010110100111", "101000110000", "111001010000", "111001010000", "001000001011", "010001101111", "011010101111", "010001101111"), 
		("010110100111", "101000110000", "111001010000", "111111111111", "001000001011", "000000010000", "010001101111", "010001101111"), 
		("010110100111", "010110100111", "101000110000", "101000110000", "001000001011", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "010110100111", "010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111")
	),
	(
		("010110100111", "010110100111", "010110100111", "010110100111", "100001000000", "100001000000", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "010110100111", "100001000000", "100001000000", "010110100111", "010110100111", "010110100111"), 
		("010110100111", "010110100111", "101000110000", "100001000000", "101000110000", "101000110000", "010110100111", "010110100111"), 
		("001000001011", "101000110000", "111111111111", "111001010000", "111001010000", "111111111111", "101000110000", "001000001011"), 
		("001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011", "001000001011"), 
		("001000001011", "010001101111", "000000010000", "010001101111", "010001101111", "000000010000", "010001101111", "001000001011"), 
		("001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "010001101111", "010001101111", "001000001011"), 
		("010110100111", "001000001011", "010001101111", "010001101111", "011010101111", "010001101111", "001000001011", "010110100111")
	),
	(
		("010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "100001000000", "010110100111", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "001000001011", "100001000000", "010110100111", "010110100111", "010110100111"), 
		("010001101111", "010001101111", "000000010000", "001000001011", "111111111111", "101000110000", "010110100111", "010110100111"), 
		("010001101111", "011010101111", "010001101111", "001000001011", "111001010000", "111001010000", "101000110000", "010110100111"), 
		("011010101111", "010001101111", "010001101111", "001000001011", "111001010000", "111001010000", "101000110000", "010110100111"), 
		("010001101111", "010001101111", "000000010000", "001000001011", "111111111111", "111001010000", "101000110000", "010110100111"), 
		("001000001011", "010001101111", "010001101111", "001000001011", "101000110000", "101000110000", "010110100111", "010110100111"), 
		("010110100111", "001000001011", "001000001011", "001000001011", "001000001011", "010110100111", "010110100111", "010110100111")
	));
begin
    data <= rom(tile_index)(to_integer(tile_offy))(to_integer(tile_offx));
end Behavioral; 